module exparser(register, result);
	input [3:0] register;
	output [3:0] result;

	assign result = register;

endmodule